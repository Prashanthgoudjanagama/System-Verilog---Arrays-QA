module PS3();



endmodule : PS2
