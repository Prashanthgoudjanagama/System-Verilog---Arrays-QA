module PS4();



endmodule : PS4
